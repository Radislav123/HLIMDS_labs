// multiprocessor_tutorial_main_system_philosopher_two.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module multiprocessor_tutorial_main_system_philosopher_two (
		output wire        cpu_jtag_debug_module_reset_reset,   // cpu_jtag_debug_module_reset.reset
		output wire        incoming_philo_slave_waitrequest,    //        incoming_philo_slave.waitrequest
		output wire [31:0] incoming_philo_slave_readdata,       //                            .readdata
		output wire        incoming_philo_slave_readdatavalid,  //                            .readdatavalid
		input  wire [0:0]  incoming_philo_slave_burstcount,     //                            .burstcount
		input  wire [31:0] incoming_philo_slave_writedata,      //                            .writedata
		input  wire [15:0] incoming_philo_slave_address,        //                            .address
		input  wire        incoming_philo_slave_write,          //                            .write
		input  wire        incoming_philo_slave_read,           //                            .read
		input  wire [3:0]  incoming_philo_slave_byteenable,     //                            .byteenable
		input  wire        incoming_philo_slave_debugaccess,    //                            .debugaccess
		input  wire        outgoing_master_waitrequest,         //             outgoing_master.waitrequest
		input  wire [31:0] outgoing_master_readdata,            //                            .readdata
		input  wire        outgoing_master_readdatavalid,       //                            .readdatavalid
		output wire [0:0]  outgoing_master_burstcount,          //                            .burstcount
		output wire [31:0] outgoing_master_writedata,           //                            .writedata
		output wire [25:0] outgoing_master_address,             //                            .address
		output wire        outgoing_master_write,               //                            .write
		output wire        outgoing_master_read,                //                            .read
		output wire [3:0]  outgoing_master_byteenable,          //                            .byteenable
		output wire        outgoing_master_debugaccess,         //                            .debugaccess
		input  wire        outgoing_philo_master_waitrequest,   //       outgoing_philo_master.waitrequest
		input  wire [31:0] outgoing_philo_master_readdata,      //                            .readdata
		input  wire        outgoing_philo_master_readdatavalid, //                            .readdatavalid
		output wire [0:0]  outgoing_philo_master_burstcount,    //                            .burstcount
		output wire [31:0] outgoing_philo_master_writedata,     //                            .writedata
		output wire [18:0] outgoing_philo_master_address,       //                            .address
		output wire        outgoing_philo_master_write,         //                            .write
		output wire        outgoing_philo_master_read,          //                            .read
		output wire [3:0]  outgoing_philo_master_byteenable,    //                            .byteenable
		output wire        outgoing_philo_master_debugaccess,   //                            .debugaccess
		input  wire        philosopher_clk_in_clk,              //          philosopher_clk_in.clk
		input  wire        philosopher_clk_reset_in_reset_n     //    philosopher_clk_reset_in.reset_n
	);

	wire  [31:0] cpu_two_data_master_readdata;                              // mm_interconnect_0:cpu_two_data_master_readdata -> cpu_two:d_readdata
	wire         cpu_two_data_master_waitrequest;                           // mm_interconnect_0:cpu_two_data_master_waitrequest -> cpu_two:d_waitrequest
	wire         cpu_two_data_master_debugaccess;                           // cpu_two:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_two_data_master_debugaccess
	wire  [26:0] cpu_two_data_master_address;                               // cpu_two:d_address -> mm_interconnect_0:cpu_two_data_master_address
	wire   [3:0] cpu_two_data_master_byteenable;                            // cpu_two:d_byteenable -> mm_interconnect_0:cpu_two_data_master_byteenable
	wire         cpu_two_data_master_read;                                  // cpu_two:d_read -> mm_interconnect_0:cpu_two_data_master_read
	wire         cpu_two_data_master_write;                                 // cpu_two:d_write -> mm_interconnect_0:cpu_two_data_master_write
	wire  [31:0] cpu_two_data_master_writedata;                             // cpu_two:d_writedata -> mm_interconnect_0:cpu_two_data_master_writedata
	wire  [31:0] cpu_two_instruction_master_readdata;                       // mm_interconnect_0:cpu_two_instruction_master_readdata -> cpu_two:i_readdata
	wire         cpu_two_instruction_master_waitrequest;                    // mm_interconnect_0:cpu_two_instruction_master_waitrequest -> cpu_two:i_waitrequest
	wire  [26:0] cpu_two_instruction_master_address;                        // cpu_two:i_address -> mm_interconnect_0:cpu_two_instruction_master_address
	wire         cpu_two_instruction_master_read;                           // cpu_two:i_read -> mm_interconnect_0:cpu_two_instruction_master_read
	wire         in_philo_bridge_m0_waitrequest;                            // mm_interconnect_0:in_philo_bridge_m0_waitrequest -> in_philo_bridge:m0_waitrequest
	wire  [31:0] in_philo_bridge_m0_readdata;                               // mm_interconnect_0:in_philo_bridge_m0_readdata -> in_philo_bridge:m0_readdata
	wire         in_philo_bridge_m0_debugaccess;                            // in_philo_bridge:m0_debugaccess -> mm_interconnect_0:in_philo_bridge_m0_debugaccess
	wire  [15:0] in_philo_bridge_m0_address;                                // in_philo_bridge:m0_address -> mm_interconnect_0:in_philo_bridge_m0_address
	wire         in_philo_bridge_m0_read;                                   // in_philo_bridge:m0_read -> mm_interconnect_0:in_philo_bridge_m0_read
	wire   [3:0] in_philo_bridge_m0_byteenable;                             // in_philo_bridge:m0_byteenable -> mm_interconnect_0:in_philo_bridge_m0_byteenable
	wire         in_philo_bridge_m0_readdatavalid;                          // mm_interconnect_0:in_philo_bridge_m0_readdatavalid -> in_philo_bridge:m0_readdatavalid
	wire  [31:0] in_philo_bridge_m0_writedata;                              // in_philo_bridge:m0_writedata -> mm_interconnect_0:in_philo_bridge_m0_writedata
	wire         in_philo_bridge_m0_write;                                  // in_philo_bridge:m0_write -> mm_interconnect_0:in_philo_bridge_m0_write
	wire   [0:0] in_philo_bridge_m0_burstcount;                             // in_philo_bridge:m0_burstcount -> mm_interconnect_0:in_philo_bridge_m0_burstcount
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_two_debug_mem_slave_readdata;        // cpu_two:debug_mem_slave_readdata -> mm_interconnect_0:cpu_two_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_two_debug_mem_slave_waitrequest;     // cpu_two:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_two_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_two_debug_mem_slave_debugaccess;     // mm_interconnect_0:cpu_two_debug_mem_slave_debugaccess -> cpu_two:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_two_debug_mem_slave_address;         // mm_interconnect_0:cpu_two_debug_mem_slave_address -> cpu_two:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_two_debug_mem_slave_read;            // mm_interconnect_0:cpu_two_debug_mem_slave_read -> cpu_two:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_two_debug_mem_slave_byteenable;      // mm_interconnect_0:cpu_two_debug_mem_slave_byteenable -> cpu_two:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_two_debug_mem_slave_write;           // mm_interconnect_0:cpu_two_debug_mem_slave_write -> cpu_two:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_two_debug_mem_slave_writedata;       // mm_interconnect_0:cpu_two_debug_mem_slave_writedata -> cpu_two:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_readdata;           // out_system_bridge:s0_readdata -> mm_interconnect_0:out_system_bridge_s0_readdata
	wire         mm_interconnect_0_out_system_bridge_s0_waitrequest;        // out_system_bridge:s0_waitrequest -> mm_interconnect_0:out_system_bridge_s0_waitrequest
	wire         mm_interconnect_0_out_system_bridge_s0_debugaccess;        // mm_interconnect_0:out_system_bridge_s0_debugaccess -> out_system_bridge:s0_debugaccess
	wire  [25:0] mm_interconnect_0_out_system_bridge_s0_address;            // mm_interconnect_0:out_system_bridge_s0_address -> out_system_bridge:s0_address
	wire         mm_interconnect_0_out_system_bridge_s0_read;               // mm_interconnect_0:out_system_bridge_s0_read -> out_system_bridge:s0_read
	wire   [3:0] mm_interconnect_0_out_system_bridge_s0_byteenable;         // mm_interconnect_0:out_system_bridge_s0_byteenable -> out_system_bridge:s0_byteenable
	wire         mm_interconnect_0_out_system_bridge_s0_readdatavalid;      // out_system_bridge:s0_readdatavalid -> mm_interconnect_0:out_system_bridge_s0_readdatavalid
	wire         mm_interconnect_0_out_system_bridge_s0_write;              // mm_interconnect_0:out_system_bridge_s0_write -> out_system_bridge:s0_write
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_writedata;          // mm_interconnect_0:out_system_bridge_s0_writedata -> out_system_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_out_system_bridge_s0_burstcount;         // mm_interconnect_0:out_system_bridge_s0_burstcount -> out_system_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_out_philo_bridge_s0_readdata;            // out_philo_bridge:s0_readdata -> mm_interconnect_0:out_philo_bridge_s0_readdata
	wire         mm_interconnect_0_out_philo_bridge_s0_waitrequest;         // out_philo_bridge:s0_waitrequest -> mm_interconnect_0:out_philo_bridge_s0_waitrequest
	wire         mm_interconnect_0_out_philo_bridge_s0_debugaccess;         // mm_interconnect_0:out_philo_bridge_s0_debugaccess -> out_philo_bridge:s0_debugaccess
	wire  [18:0] mm_interconnect_0_out_philo_bridge_s0_address;             // mm_interconnect_0:out_philo_bridge_s0_address -> out_philo_bridge:s0_address
	wire         mm_interconnect_0_out_philo_bridge_s0_read;                // mm_interconnect_0:out_philo_bridge_s0_read -> out_philo_bridge:s0_read
	wire   [3:0] mm_interconnect_0_out_philo_bridge_s0_byteenable;          // mm_interconnect_0:out_philo_bridge_s0_byteenable -> out_philo_bridge:s0_byteenable
	wire         mm_interconnect_0_out_philo_bridge_s0_readdatavalid;       // out_philo_bridge:s0_readdatavalid -> mm_interconnect_0:out_philo_bridge_s0_readdatavalid
	wire         mm_interconnect_0_out_philo_bridge_s0_write;               // mm_interconnect_0:out_philo_bridge_s0_write -> out_philo_bridge:s0_write
	wire  [31:0] mm_interconnect_0_out_philo_bridge_s0_writedata;           // mm_interconnect_0:out_philo_bridge_s0_writedata -> out_philo_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_out_philo_bridge_s0_burstcount;          // mm_interconnect_0:out_philo_bridge_s0_burstcount -> out_philo_bridge:s0_burstcount
	wire         mm_interconnect_0_chopstick_mutex_s1_chipselect;           // mm_interconnect_0:chopstick_mutex_s1_chipselect -> chopstick_mutex:chipselect
	wire  [31:0] mm_interconnect_0_chopstick_mutex_s1_readdata;             // chopstick_mutex:data_to_cpu -> mm_interconnect_0:chopstick_mutex_s1_readdata
	wire   [0:0] mm_interconnect_0_chopstick_mutex_s1_address;              // mm_interconnect_0:chopstick_mutex_s1_address -> chopstick_mutex:address
	wire         mm_interconnect_0_chopstick_mutex_s1_read;                 // mm_interconnect_0:chopstick_mutex_s1_read -> chopstick_mutex:read
	wire         mm_interconnect_0_chopstick_mutex_s1_write;                // mm_interconnect_0:chopstick_mutex_s1_write -> chopstick_mutex:write
	wire  [31:0] mm_interconnect_0_chopstick_mutex_s1_writedata;            // mm_interconnect_0:chopstick_mutex_s1_writedata -> chopstick_mutex:data_from_cpu
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         irq_mapper_receiver0_irq;                                  // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_two_irq_irq;                                           // irq_mapper:sender_irq -> cpu_two:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [chopstick_mutex:reset_n, cpu_two:reset_n, in_philo_bridge:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_two_reset_reset_bridge_in_reset_reset, out_philo_bridge:reset, out_system_bridge:reset, rst_translator:in_reset, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu_two:reset_req, rst_translator:reset_req_in]

	multiprocessor_tutorial_main_system_philosopher_one_chopstick_mutex chopstick_mutex (
		.reset_n       (~rst_controller_reset_out_reset),                 // reset.reset_n
		.clk           (philosopher_clk_in_clk),                          //   clk.clk
		.chipselect    (mm_interconnect_0_chopstick_mutex_s1_chipselect), //    s1.chipselect
		.data_from_cpu (mm_interconnect_0_chopstick_mutex_s1_writedata),  //      .writedata
		.read          (mm_interconnect_0_chopstick_mutex_s1_read),       //      .read
		.write         (mm_interconnect_0_chopstick_mutex_s1_write),      //      .write
		.data_to_cpu   (mm_interconnect_0_chopstick_mutex_s1_readdata),   //      .readdata
		.address       (mm_interconnect_0_chopstick_mutex_s1_address)     //      .address
	);

	multiprocessor_tutorial_main_system_philosopher_two_cpu_two cpu_two (
		.clk                                 (philosopher_clk_in_clk),                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (cpu_two_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_two_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_two_data_master_read),                              //                          .read
		.d_readdata                          (cpu_two_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_two_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_two_data_master_write),                             //                          .write
		.d_writedata                         (cpu_two_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_two_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_two_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_two_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_two_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_two_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_two_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_jtag_debug_module_reset_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_two_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_two_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_two_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_two_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_two_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_two_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_two_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_two_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (16),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) in_philo_bridge (
		.clk              (philosopher_clk_in_clk),             //   clk.clk
		.reset            (rst_controller_reset_out_reset),     // reset.reset
		.s0_waitrequest   (incoming_philo_slave_waitrequest),   //    s0.waitrequest
		.s0_readdata      (incoming_philo_slave_readdata),      //      .readdata
		.s0_readdatavalid (incoming_philo_slave_readdatavalid), //      .readdatavalid
		.s0_burstcount    (incoming_philo_slave_burstcount),    //      .burstcount
		.s0_writedata     (incoming_philo_slave_writedata),     //      .writedata
		.s0_address       (incoming_philo_slave_address),       //      .address
		.s0_write         (incoming_philo_slave_write),         //      .write
		.s0_read          (incoming_philo_slave_read),          //      .read
		.s0_byteenable    (incoming_philo_slave_byteenable),    //      .byteenable
		.s0_debugaccess   (incoming_philo_slave_debugaccess),   //      .debugaccess
		.m0_waitrequest   (in_philo_bridge_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (in_philo_bridge_m0_readdata),        //      .readdata
		.m0_readdatavalid (in_philo_bridge_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (in_philo_bridge_m0_burstcount),      //      .burstcount
		.m0_writedata     (in_philo_bridge_m0_writedata),       //      .writedata
		.m0_address       (in_philo_bridge_m0_address),         //      .address
		.m0_write         (in_philo_bridge_m0_write),           //      .write
		.m0_read          (in_philo_bridge_m0_read),            //      .read
		.m0_byteenable    (in_philo_bridge_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (in_philo_bridge_m0_debugaccess),     //      .debugaccess
		.s0_response      (),                                   // (terminated)
		.m0_response      (2'b00)                               // (terminated)
	);

	multiprocessor_tutorial_main_system_jtag_uart_top jtag_uart (
		.clk            (philosopher_clk_in_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (19),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) out_philo_bridge (
		.clk              (philosopher_clk_in_clk),                              //   clk.clk
		.reset            (rst_controller_reset_out_reset),                      // reset.reset
		.s0_waitrequest   (mm_interconnect_0_out_philo_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_out_philo_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_out_philo_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_out_philo_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_out_philo_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_out_philo_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_out_philo_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_out_philo_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_out_philo_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_out_philo_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (outgoing_philo_master_waitrequest),                   //    m0.waitrequest
		.m0_readdata      (outgoing_philo_master_readdata),                      //      .readdata
		.m0_readdatavalid (outgoing_philo_master_readdatavalid),                 //      .readdatavalid
		.m0_burstcount    (outgoing_philo_master_burstcount),                    //      .burstcount
		.m0_writedata     (outgoing_philo_master_writedata),                     //      .writedata
		.m0_address       (outgoing_philo_master_address),                       //      .address
		.m0_write         (outgoing_philo_master_write),                         //      .write
		.m0_read          (outgoing_philo_master_read),                          //      .read
		.m0_byteenable    (outgoing_philo_master_byteenable),                    //      .byteenable
		.m0_debugaccess   (outgoing_philo_master_debugaccess),                   //      .debugaccess
		.s0_response      (),                                                    // (terminated)
		.m0_response      (2'b00)                                                // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (26),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) out_system_bridge (
		.clk              (philosopher_clk_in_clk),                               //   clk.clk
		.reset            (rst_controller_reset_out_reset),                       // reset.reset
		.s0_waitrequest   (mm_interconnect_0_out_system_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_out_system_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_out_system_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_out_system_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_out_system_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_out_system_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_out_system_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_out_system_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_out_system_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_out_system_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (outgoing_master_waitrequest),                          //    m0.waitrequest
		.m0_readdata      (outgoing_master_readdata),                             //      .readdata
		.m0_readdatavalid (outgoing_master_readdatavalid),                        //      .readdatavalid
		.m0_burstcount    (outgoing_master_burstcount),                           //      .burstcount
		.m0_writedata     (outgoing_master_writedata),                            //      .writedata
		.m0_address       (outgoing_master_address),                              //      .address
		.m0_write         (outgoing_master_write),                                //      .write
		.m0_read          (outgoing_master_read),                                 //      .read
		.m0_byteenable    (outgoing_master_byteenable),                           //      .byteenable
		.m0_debugaccess   (outgoing_master_debugaccess),                          //      .debugaccess
		.s0_response      (),                                                     // (terminated)
		.m0_response      (2'b00)                                                 // (terminated)
	);

	multiprocessor_tutorial_main_system_timer_top timer (
		.clk        (philosopher_clk_in_clk),                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	multiprocessor_tutorial_main_system_philosopher_two_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                               (philosopher_clk_in_clk),                                    //                             clk_clk.clk
		.cpu_two_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpu_two_reset_reset_bridge_in_reset.reset
		.cpu_two_data_master_address               (cpu_two_data_master_address),                               //                 cpu_two_data_master.address
		.cpu_two_data_master_waitrequest           (cpu_two_data_master_waitrequest),                           //                                    .waitrequest
		.cpu_two_data_master_byteenable            (cpu_two_data_master_byteenable),                            //                                    .byteenable
		.cpu_two_data_master_read                  (cpu_two_data_master_read),                                  //                                    .read
		.cpu_two_data_master_readdata              (cpu_two_data_master_readdata),                              //                                    .readdata
		.cpu_two_data_master_write                 (cpu_two_data_master_write),                                 //                                    .write
		.cpu_two_data_master_writedata             (cpu_two_data_master_writedata),                             //                                    .writedata
		.cpu_two_data_master_debugaccess           (cpu_two_data_master_debugaccess),                           //                                    .debugaccess
		.cpu_two_instruction_master_address        (cpu_two_instruction_master_address),                        //          cpu_two_instruction_master.address
		.cpu_two_instruction_master_waitrequest    (cpu_two_instruction_master_waitrequest),                    //                                    .waitrequest
		.cpu_two_instruction_master_read           (cpu_two_instruction_master_read),                           //                                    .read
		.cpu_two_instruction_master_readdata       (cpu_two_instruction_master_readdata),                       //                                    .readdata
		.in_philo_bridge_m0_address                (in_philo_bridge_m0_address),                                //                  in_philo_bridge_m0.address
		.in_philo_bridge_m0_waitrequest            (in_philo_bridge_m0_waitrequest),                            //                                    .waitrequest
		.in_philo_bridge_m0_burstcount             (in_philo_bridge_m0_burstcount),                             //                                    .burstcount
		.in_philo_bridge_m0_byteenable             (in_philo_bridge_m0_byteenable),                             //                                    .byteenable
		.in_philo_bridge_m0_read                   (in_philo_bridge_m0_read),                                   //                                    .read
		.in_philo_bridge_m0_readdata               (in_philo_bridge_m0_readdata),                               //                                    .readdata
		.in_philo_bridge_m0_readdatavalid          (in_philo_bridge_m0_readdatavalid),                          //                                    .readdatavalid
		.in_philo_bridge_m0_write                  (in_philo_bridge_m0_write),                                  //                                    .write
		.in_philo_bridge_m0_writedata              (in_philo_bridge_m0_writedata),                              //                                    .writedata
		.in_philo_bridge_m0_debugaccess            (in_philo_bridge_m0_debugaccess),                            //                                    .debugaccess
		.chopstick_mutex_s1_address                (mm_interconnect_0_chopstick_mutex_s1_address),              //                  chopstick_mutex_s1.address
		.chopstick_mutex_s1_write                  (mm_interconnect_0_chopstick_mutex_s1_write),                //                                    .write
		.chopstick_mutex_s1_read                   (mm_interconnect_0_chopstick_mutex_s1_read),                 //                                    .read
		.chopstick_mutex_s1_readdata               (mm_interconnect_0_chopstick_mutex_s1_readdata),             //                                    .readdata
		.chopstick_mutex_s1_writedata              (mm_interconnect_0_chopstick_mutex_s1_writedata),            //                                    .writedata
		.chopstick_mutex_s1_chipselect             (mm_interconnect_0_chopstick_mutex_s1_chipselect),           //                                    .chipselect
		.cpu_two_debug_mem_slave_address           (mm_interconnect_0_cpu_two_debug_mem_slave_address),         //             cpu_two_debug_mem_slave.address
		.cpu_two_debug_mem_slave_write             (mm_interconnect_0_cpu_two_debug_mem_slave_write),           //                                    .write
		.cpu_two_debug_mem_slave_read              (mm_interconnect_0_cpu_two_debug_mem_slave_read),            //                                    .read
		.cpu_two_debug_mem_slave_readdata          (mm_interconnect_0_cpu_two_debug_mem_slave_readdata),        //                                    .readdata
		.cpu_two_debug_mem_slave_writedata         (mm_interconnect_0_cpu_two_debug_mem_slave_writedata),       //                                    .writedata
		.cpu_two_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_two_debug_mem_slave_byteenable),      //                                    .byteenable
		.cpu_two_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_two_debug_mem_slave_waitrequest),     //                                    .waitrequest
		.cpu_two_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_two_debug_mem_slave_debugaccess),     //                                    .debugaccess
		.jtag_uart_avalon_jtag_slave_address       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                    .write
		.jtag_uart_avalon_jtag_slave_read          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                    .read
		.jtag_uart_avalon_jtag_slave_readdata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.out_philo_bridge_s0_address               (mm_interconnect_0_out_philo_bridge_s0_address),             //                 out_philo_bridge_s0.address
		.out_philo_bridge_s0_write                 (mm_interconnect_0_out_philo_bridge_s0_write),               //                                    .write
		.out_philo_bridge_s0_read                  (mm_interconnect_0_out_philo_bridge_s0_read),                //                                    .read
		.out_philo_bridge_s0_readdata              (mm_interconnect_0_out_philo_bridge_s0_readdata),            //                                    .readdata
		.out_philo_bridge_s0_writedata             (mm_interconnect_0_out_philo_bridge_s0_writedata),           //                                    .writedata
		.out_philo_bridge_s0_burstcount            (mm_interconnect_0_out_philo_bridge_s0_burstcount),          //                                    .burstcount
		.out_philo_bridge_s0_byteenable            (mm_interconnect_0_out_philo_bridge_s0_byteenable),          //                                    .byteenable
		.out_philo_bridge_s0_readdatavalid         (mm_interconnect_0_out_philo_bridge_s0_readdatavalid),       //                                    .readdatavalid
		.out_philo_bridge_s0_waitrequest           (mm_interconnect_0_out_philo_bridge_s0_waitrequest),         //                                    .waitrequest
		.out_philo_bridge_s0_debugaccess           (mm_interconnect_0_out_philo_bridge_s0_debugaccess),         //                                    .debugaccess
		.out_system_bridge_s0_address              (mm_interconnect_0_out_system_bridge_s0_address),            //                out_system_bridge_s0.address
		.out_system_bridge_s0_write                (mm_interconnect_0_out_system_bridge_s0_write),              //                                    .write
		.out_system_bridge_s0_read                 (mm_interconnect_0_out_system_bridge_s0_read),               //                                    .read
		.out_system_bridge_s0_readdata             (mm_interconnect_0_out_system_bridge_s0_readdata),           //                                    .readdata
		.out_system_bridge_s0_writedata            (mm_interconnect_0_out_system_bridge_s0_writedata),          //                                    .writedata
		.out_system_bridge_s0_burstcount           (mm_interconnect_0_out_system_bridge_s0_burstcount),         //                                    .burstcount
		.out_system_bridge_s0_byteenable           (mm_interconnect_0_out_system_bridge_s0_byteenable),         //                                    .byteenable
		.out_system_bridge_s0_readdatavalid        (mm_interconnect_0_out_system_bridge_s0_readdatavalid),      //                                    .readdatavalid
		.out_system_bridge_s0_waitrequest          (mm_interconnect_0_out_system_bridge_s0_waitrequest),        //                                    .waitrequest
		.out_system_bridge_s0_debugaccess          (mm_interconnect_0_out_system_bridge_s0_debugaccess),        //                                    .debugaccess
		.timer_s1_address                          (mm_interconnect_0_timer_s1_address),                        //                            timer_s1.address
		.timer_s1_write                            (mm_interconnect_0_timer_s1_write),                          //                                    .write
		.timer_s1_readdata                         (mm_interconnect_0_timer_s1_readdata),                       //                                    .readdata
		.timer_s1_writedata                        (mm_interconnect_0_timer_s1_writedata),                      //                                    .writedata
		.timer_s1_chipselect                       (mm_interconnect_0_timer_s1_chipselect)                      //                                    .chipselect
	);

	multiprocessor_tutorial_main_system_irq_mapper irq_mapper (
		.clk           (philosopher_clk_in_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_two_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~philosopher_clk_reset_in_reset_n),  // reset_in0.reset
		.clk            (philosopher_clk_in_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
