
module multiprocessor_tutorial_main_system (
	clk_clk_in_reset_reset_n,
	clk_in_clk);	

	input		clk_clk_in_reset_reset_n;
	input		clk_in_clk;
endmodule
