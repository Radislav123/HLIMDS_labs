// multiprocessor_tutorial_main_system.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module multiprocessor_tutorial_main_system (
		input  wire  clk_clk_in_reset_reset_n, // clk_clk_in_reset.reset_n
		input  wire  clk_in_clk                //           clk_in.clk
	);

	wire  [31:0] cpu_top_data_master_readdata;                                          // mm_interconnect_0:cpu_top_data_master_readdata -> cpu_top:d_readdata
	wire         cpu_top_data_master_waitrequest;                                       // mm_interconnect_0:cpu_top_data_master_waitrequest -> cpu_top:d_waitrequest
	wire         cpu_top_data_master_debugaccess;                                       // cpu_top:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_top_data_master_debugaccess
	wire  [18:0] cpu_top_data_master_address;                                           // cpu_top:d_address -> mm_interconnect_0:cpu_top_data_master_address
	wire   [3:0] cpu_top_data_master_byteenable;                                        // cpu_top:d_byteenable -> mm_interconnect_0:cpu_top_data_master_byteenable
	wire         cpu_top_data_master_read;                                              // cpu_top:d_read -> mm_interconnect_0:cpu_top_data_master_read
	wire         cpu_top_data_master_write;                                             // cpu_top:d_write -> mm_interconnect_0:cpu_top_data_master_write
	wire  [31:0] cpu_top_data_master_writedata;                                         // cpu_top:d_writedata -> mm_interconnect_0:cpu_top_data_master_writedata
	wire  [31:0] cpu_top_instruction_master_readdata;                                   // mm_interconnect_0:cpu_top_instruction_master_readdata -> cpu_top:i_readdata
	wire         cpu_top_instruction_master_waitrequest;                                // mm_interconnect_0:cpu_top_instruction_master_waitrequest -> cpu_top:i_waitrequest
	wire  [18:0] cpu_top_instruction_master_address;                                    // cpu_top:i_address -> mm_interconnect_0:cpu_top_instruction_master_address
	wire         cpu_top_instruction_master_read;                                       // cpu_top:i_read -> mm_interconnect_0:cpu_top_instruction_master_read
	wire         philosopher_two_outgoing_master_waitrequest;                           // mm_interconnect_0:philosopher_two_outgoing_master_waitrequest -> philosopher_two:outgoing_master_waitrequest
	wire  [31:0] philosopher_two_outgoing_master_readdata;                              // mm_interconnect_0:philosopher_two_outgoing_master_readdata -> philosopher_two:outgoing_master_readdata
	wire         philosopher_two_outgoing_master_debugaccess;                           // philosopher_two:outgoing_master_debugaccess -> mm_interconnect_0:philosopher_two_outgoing_master_debugaccess
	wire  [25:0] philosopher_two_outgoing_master_address;                               // philosopher_two:outgoing_master_address -> mm_interconnect_0:philosopher_two_outgoing_master_address
	wire         philosopher_two_outgoing_master_read;                                  // philosopher_two:outgoing_master_read -> mm_interconnect_0:philosopher_two_outgoing_master_read
	wire   [3:0] philosopher_two_outgoing_master_byteenable;                            // philosopher_two:outgoing_master_byteenable -> mm_interconnect_0:philosopher_two_outgoing_master_byteenable
	wire         philosopher_two_outgoing_master_readdatavalid;                         // mm_interconnect_0:philosopher_two_outgoing_master_readdatavalid -> philosopher_two:outgoing_master_readdatavalid
	wire  [31:0] philosopher_two_outgoing_master_writedata;                             // philosopher_two:outgoing_master_writedata -> mm_interconnect_0:philosopher_two_outgoing_master_writedata
	wire         philosopher_two_outgoing_master_write;                                 // philosopher_two:outgoing_master_write -> mm_interconnect_0:philosopher_two_outgoing_master_write
	wire   [0:0] philosopher_two_outgoing_master_burstcount;                            // philosopher_two:outgoing_master_burstcount -> mm_interconnect_0:philosopher_two_outgoing_master_burstcount
	wire         philosopher_one_outgoing_master_waitrequest;                           // mm_interconnect_0:philosopher_one_outgoing_master_waitrequest -> philosopher_one:outgoing_master_waitrequest
	wire  [31:0] philosopher_one_outgoing_master_readdata;                              // mm_interconnect_0:philosopher_one_outgoing_master_readdata -> philosopher_one:outgoing_master_readdata
	wire         philosopher_one_outgoing_master_debugaccess;                           // philosopher_one:outgoing_master_debugaccess -> mm_interconnect_0:philosopher_one_outgoing_master_debugaccess
	wire  [25:0] philosopher_one_outgoing_master_address;                               // philosopher_one:outgoing_master_address -> mm_interconnect_0:philosopher_one_outgoing_master_address
	wire         philosopher_one_outgoing_master_read;                                  // philosopher_one:outgoing_master_read -> mm_interconnect_0:philosopher_one_outgoing_master_read
	wire   [3:0] philosopher_one_outgoing_master_byteenable;                            // philosopher_one:outgoing_master_byteenable -> mm_interconnect_0:philosopher_one_outgoing_master_byteenable
	wire         philosopher_one_outgoing_master_readdatavalid;                         // mm_interconnect_0:philosopher_one_outgoing_master_readdatavalid -> philosopher_one:outgoing_master_readdatavalid
	wire  [31:0] philosopher_one_outgoing_master_writedata;                             // philosopher_one:outgoing_master_writedata -> mm_interconnect_0:philosopher_one_outgoing_master_writedata
	wire         philosopher_one_outgoing_master_write;                                 // philosopher_one:outgoing_master_write -> mm_interconnect_0:philosopher_one_outgoing_master_write
	wire   [0:0] philosopher_one_outgoing_master_burstcount;                            // philosopher_one:outgoing_master_burstcount -> mm_interconnect_0:philosopher_one_outgoing_master_burstcount
	wire         philosopher_zero_outgoing_master_waitrequest;                          // mm_interconnect_0:philosopher_zero_outgoing_master_waitrequest -> philosopher_zero:outgoing_master_waitrequest
	wire  [31:0] philosopher_zero_outgoing_master_readdata;                             // mm_interconnect_0:philosopher_zero_outgoing_master_readdata -> philosopher_zero:outgoing_master_readdata
	wire         philosopher_zero_outgoing_master_debugaccess;                          // philosopher_zero:outgoing_master_debugaccess -> mm_interconnect_0:philosopher_zero_outgoing_master_debugaccess
	wire  [25:0] philosopher_zero_outgoing_master_address;                              // philosopher_zero:outgoing_master_address -> mm_interconnect_0:philosopher_zero_outgoing_master_address
	wire         philosopher_zero_outgoing_master_read;                                 // philosopher_zero:outgoing_master_read -> mm_interconnect_0:philosopher_zero_outgoing_master_read
	wire   [3:0] philosopher_zero_outgoing_master_byteenable;                           // philosopher_zero:outgoing_master_byteenable -> mm_interconnect_0:philosopher_zero_outgoing_master_byteenable
	wire         philosopher_zero_outgoing_master_readdatavalid;                        // mm_interconnect_0:philosopher_zero_outgoing_master_readdatavalid -> philosopher_zero:outgoing_master_readdatavalid
	wire  [31:0] philosopher_zero_outgoing_master_writedata;                            // philosopher_zero:outgoing_master_writedata -> mm_interconnect_0:philosopher_zero_outgoing_master_writedata
	wire         philosopher_zero_outgoing_master_write;                                // philosopher_zero:outgoing_master_write -> mm_interconnect_0:philosopher_zero_outgoing_master_write
	wire   [0:0] philosopher_zero_outgoing_master_burstcount;                           // philosopher_zero:outgoing_master_burstcount -> mm_interconnect_0:philosopher_zero_outgoing_master_burstcount
	wire         philosopher_one_outgoing_philo_master_waitrequest;                     // mm_interconnect_0:philosopher_one_outgoing_philo_master_waitrequest -> philosopher_one:outgoing_philo_master_waitrequest
	wire  [31:0] philosopher_one_outgoing_philo_master_readdata;                        // mm_interconnect_0:philosopher_one_outgoing_philo_master_readdata -> philosopher_one:outgoing_philo_master_readdata
	wire         philosopher_one_outgoing_philo_master_debugaccess;                     // philosopher_one:outgoing_philo_master_debugaccess -> mm_interconnect_0:philosopher_one_outgoing_philo_master_debugaccess
	wire  [18:0] philosopher_one_outgoing_philo_master_address;                         // philosopher_one:outgoing_philo_master_address -> mm_interconnect_0:philosopher_one_outgoing_philo_master_address
	wire         philosopher_one_outgoing_philo_master_read;                            // philosopher_one:outgoing_philo_master_read -> mm_interconnect_0:philosopher_one_outgoing_philo_master_read
	wire   [3:0] philosopher_one_outgoing_philo_master_byteenable;                      // philosopher_one:outgoing_philo_master_byteenable -> mm_interconnect_0:philosopher_one_outgoing_philo_master_byteenable
	wire         philosopher_one_outgoing_philo_master_readdatavalid;                   // mm_interconnect_0:philosopher_one_outgoing_philo_master_readdatavalid -> philosopher_one:outgoing_philo_master_readdatavalid
	wire  [31:0] philosopher_one_outgoing_philo_master_writedata;                       // philosopher_one:outgoing_philo_master_writedata -> mm_interconnect_0:philosopher_one_outgoing_philo_master_writedata
	wire         philosopher_one_outgoing_philo_master_write;                           // philosopher_one:outgoing_philo_master_write -> mm_interconnect_0:philosopher_one_outgoing_philo_master_write
	wire   [0:0] philosopher_one_outgoing_philo_master_burstcount;                      // philosopher_one:outgoing_philo_master_burstcount -> mm_interconnect_0:philosopher_one_outgoing_philo_master_burstcount
	wire         philosopher_zero_outgoing_philo_master_waitrequest;                    // mm_interconnect_0:philosopher_zero_outgoing_philo_master_waitrequest -> philosopher_zero:outgoing_philo_master_waitrequest
	wire  [31:0] philosopher_zero_outgoing_philo_master_readdata;                       // mm_interconnect_0:philosopher_zero_outgoing_philo_master_readdata -> philosopher_zero:outgoing_philo_master_readdata
	wire         philosopher_zero_outgoing_philo_master_debugaccess;                    // philosopher_zero:outgoing_philo_master_debugaccess -> mm_interconnect_0:philosopher_zero_outgoing_philo_master_debugaccess
	wire  [18:0] philosopher_zero_outgoing_philo_master_address;                        // philosopher_zero:outgoing_philo_master_address -> mm_interconnect_0:philosopher_zero_outgoing_philo_master_address
	wire         philosopher_zero_outgoing_philo_master_read;                           // philosopher_zero:outgoing_philo_master_read -> mm_interconnect_0:philosopher_zero_outgoing_philo_master_read
	wire   [3:0] philosopher_zero_outgoing_philo_master_byteenable;                     // philosopher_zero:outgoing_philo_master_byteenable -> mm_interconnect_0:philosopher_zero_outgoing_philo_master_byteenable
	wire         philosopher_zero_outgoing_philo_master_readdatavalid;                  // mm_interconnect_0:philosopher_zero_outgoing_philo_master_readdatavalid -> philosopher_zero:outgoing_philo_master_readdatavalid
	wire  [31:0] philosopher_zero_outgoing_philo_master_writedata;                      // philosopher_zero:outgoing_philo_master_writedata -> mm_interconnect_0:philosopher_zero_outgoing_philo_master_writedata
	wire         philosopher_zero_outgoing_philo_master_write;                          // philosopher_zero:outgoing_philo_master_write -> mm_interconnect_0:philosopher_zero_outgoing_philo_master_write
	wire   [0:0] philosopher_zero_outgoing_philo_master_burstcount;                     // philosopher_zero:outgoing_philo_master_burstcount -> mm_interconnect_0:philosopher_zero_outgoing_philo_master_burstcount
	wire         philosopher_two_outgoing_philo_master_waitrequest;                     // mm_interconnect_0:philosopher_two_outgoing_philo_master_waitrequest -> philosopher_two:outgoing_philo_master_waitrequest
	wire  [31:0] philosopher_two_outgoing_philo_master_readdata;                        // mm_interconnect_0:philosopher_two_outgoing_philo_master_readdata -> philosopher_two:outgoing_philo_master_readdata
	wire         philosopher_two_outgoing_philo_master_debugaccess;                     // philosopher_two:outgoing_philo_master_debugaccess -> mm_interconnect_0:philosopher_two_outgoing_philo_master_debugaccess
	wire  [18:0] philosopher_two_outgoing_philo_master_address;                         // philosopher_two:outgoing_philo_master_address -> mm_interconnect_0:philosopher_two_outgoing_philo_master_address
	wire         philosopher_two_outgoing_philo_master_read;                            // philosopher_two:outgoing_philo_master_read -> mm_interconnect_0:philosopher_two_outgoing_philo_master_read
	wire   [3:0] philosopher_two_outgoing_philo_master_byteenable;                      // philosopher_two:outgoing_philo_master_byteenable -> mm_interconnect_0:philosopher_two_outgoing_philo_master_byteenable
	wire         philosopher_two_outgoing_philo_master_readdatavalid;                   // mm_interconnect_0:philosopher_two_outgoing_philo_master_readdatavalid -> philosopher_two:outgoing_philo_master_readdatavalid
	wire  [31:0] philosopher_two_outgoing_philo_master_writedata;                       // philosopher_two:outgoing_philo_master_writedata -> mm_interconnect_0:philosopher_two_outgoing_philo_master_writedata
	wire         philosopher_two_outgoing_philo_master_write;                           // philosopher_two:outgoing_philo_master_write -> mm_interconnect_0:philosopher_two_outgoing_philo_master_write
	wire   [0:0] philosopher_two_outgoing_philo_master_burstcount;                      // philosopher_two:outgoing_philo_master_burstcount -> mm_interconnect_0:philosopher_two_outgoing_philo_master_burstcount
	wire         mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_top_avalon_jtag_slave_chipselect -> jtag_uart_top:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_readdata;            // jtag_uart_top:av_readdata -> mm_interconnect_0:jtag_uart_top_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_waitrequest;         // jtag_uart_top:av_waitrequest -> mm_interconnect_0:jtag_uart_top_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_top_avalon_jtag_slave_address -> jtag_uart_top:av_address
	wire         mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_top_avalon_jtag_slave_read -> jtag_uart_top:av_read_n
	wire         mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_top_avalon_jtag_slave_write -> jtag_uart_top:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_top_avalon_jtag_slave_writedata -> jtag_uart_top:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                   // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                    // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_cpu_top_debug_mem_slave_readdata;                    // cpu_top:debug_mem_slave_readdata -> mm_interconnect_0:cpu_top_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_top_debug_mem_slave_waitrequest;                 // cpu_top:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_top_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_top_debug_mem_slave_debugaccess;                 // mm_interconnect_0:cpu_top_debug_mem_slave_debugaccess -> cpu_top:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_top_debug_mem_slave_address;                     // mm_interconnect_0:cpu_top_debug_mem_slave_address -> cpu_top:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_top_debug_mem_slave_read;                        // mm_interconnect_0:cpu_top_debug_mem_slave_read -> cpu_top:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_top_debug_mem_slave_byteenable;                  // mm_interconnect_0:cpu_top_debug_mem_slave_byteenable -> cpu_top:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_top_debug_mem_slave_write;                       // mm_interconnect_0:cpu_top_debug_mem_slave_write -> cpu_top:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_top_debug_mem_slave_writedata;                   // mm_interconnect_0:cpu_top_debug_mem_slave_writedata -> cpu_top:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_philosopher_zero_incoming_philo_slave_readdata;      // philosopher_zero:incoming_philo_slave_readdata -> mm_interconnect_0:philosopher_zero_incoming_philo_slave_readdata
	wire         mm_interconnect_0_philosopher_zero_incoming_philo_slave_waitrequest;   // philosopher_zero:incoming_philo_slave_waitrequest -> mm_interconnect_0:philosopher_zero_incoming_philo_slave_waitrequest
	wire         mm_interconnect_0_philosopher_zero_incoming_philo_slave_debugaccess;   // mm_interconnect_0:philosopher_zero_incoming_philo_slave_debugaccess -> philosopher_zero:incoming_philo_slave_debugaccess
	wire  [15:0] mm_interconnect_0_philosopher_zero_incoming_philo_slave_address;       // mm_interconnect_0:philosopher_zero_incoming_philo_slave_address -> philosopher_zero:incoming_philo_slave_address
	wire         mm_interconnect_0_philosopher_zero_incoming_philo_slave_read;          // mm_interconnect_0:philosopher_zero_incoming_philo_slave_read -> philosopher_zero:incoming_philo_slave_read
	wire   [3:0] mm_interconnect_0_philosopher_zero_incoming_philo_slave_byteenable;    // mm_interconnect_0:philosopher_zero_incoming_philo_slave_byteenable -> philosopher_zero:incoming_philo_slave_byteenable
	wire         mm_interconnect_0_philosopher_zero_incoming_philo_slave_readdatavalid; // philosopher_zero:incoming_philo_slave_readdatavalid -> mm_interconnect_0:philosopher_zero_incoming_philo_slave_readdatavalid
	wire         mm_interconnect_0_philosopher_zero_incoming_philo_slave_write;         // mm_interconnect_0:philosopher_zero_incoming_philo_slave_write -> philosopher_zero:incoming_philo_slave_write
	wire  [31:0] mm_interconnect_0_philosopher_zero_incoming_philo_slave_writedata;     // mm_interconnect_0:philosopher_zero_incoming_philo_slave_writedata -> philosopher_zero:incoming_philo_slave_writedata
	wire   [0:0] mm_interconnect_0_philosopher_zero_incoming_philo_slave_burstcount;    // mm_interconnect_0:philosopher_zero_incoming_philo_slave_burstcount -> philosopher_zero:incoming_philo_slave_burstcount
	wire  [31:0] mm_interconnect_0_philosopher_one_incoming_philo_slave_readdata;       // philosopher_one:incoming_philo_slave_readdata -> mm_interconnect_0:philosopher_one_incoming_philo_slave_readdata
	wire         mm_interconnect_0_philosopher_one_incoming_philo_slave_waitrequest;    // philosopher_one:incoming_philo_slave_waitrequest -> mm_interconnect_0:philosopher_one_incoming_philo_slave_waitrequest
	wire         mm_interconnect_0_philosopher_one_incoming_philo_slave_debugaccess;    // mm_interconnect_0:philosopher_one_incoming_philo_slave_debugaccess -> philosopher_one:incoming_philo_slave_debugaccess
	wire  [15:0] mm_interconnect_0_philosopher_one_incoming_philo_slave_address;        // mm_interconnect_0:philosopher_one_incoming_philo_slave_address -> philosopher_one:incoming_philo_slave_address
	wire         mm_interconnect_0_philosopher_one_incoming_philo_slave_read;           // mm_interconnect_0:philosopher_one_incoming_philo_slave_read -> philosopher_one:incoming_philo_slave_read
	wire   [3:0] mm_interconnect_0_philosopher_one_incoming_philo_slave_byteenable;     // mm_interconnect_0:philosopher_one_incoming_philo_slave_byteenable -> philosopher_one:incoming_philo_slave_byteenable
	wire         mm_interconnect_0_philosopher_one_incoming_philo_slave_readdatavalid;  // philosopher_one:incoming_philo_slave_readdatavalid -> mm_interconnect_0:philosopher_one_incoming_philo_slave_readdatavalid
	wire         mm_interconnect_0_philosopher_one_incoming_philo_slave_write;          // mm_interconnect_0:philosopher_one_incoming_philo_slave_write -> philosopher_one:incoming_philo_slave_write
	wire  [31:0] mm_interconnect_0_philosopher_one_incoming_philo_slave_writedata;      // mm_interconnect_0:philosopher_one_incoming_philo_slave_writedata -> philosopher_one:incoming_philo_slave_writedata
	wire   [0:0] mm_interconnect_0_philosopher_one_incoming_philo_slave_burstcount;     // mm_interconnect_0:philosopher_one_incoming_philo_slave_burstcount -> philosopher_one:incoming_philo_slave_burstcount
	wire  [31:0] mm_interconnect_0_philosopher_two_incoming_philo_slave_readdata;       // philosopher_two:incoming_philo_slave_readdata -> mm_interconnect_0:philosopher_two_incoming_philo_slave_readdata
	wire         mm_interconnect_0_philosopher_two_incoming_philo_slave_waitrequest;    // philosopher_two:incoming_philo_slave_waitrequest -> mm_interconnect_0:philosopher_two_incoming_philo_slave_waitrequest
	wire         mm_interconnect_0_philosopher_two_incoming_philo_slave_debugaccess;    // mm_interconnect_0:philosopher_two_incoming_philo_slave_debugaccess -> philosopher_two:incoming_philo_slave_debugaccess
	wire  [15:0] mm_interconnect_0_philosopher_two_incoming_philo_slave_address;        // mm_interconnect_0:philosopher_two_incoming_philo_slave_address -> philosopher_two:incoming_philo_slave_address
	wire         mm_interconnect_0_philosopher_two_incoming_philo_slave_read;           // mm_interconnect_0:philosopher_two_incoming_philo_slave_read -> philosopher_two:incoming_philo_slave_read
	wire   [3:0] mm_interconnect_0_philosopher_two_incoming_philo_slave_byteenable;     // mm_interconnect_0:philosopher_two_incoming_philo_slave_byteenable -> philosopher_two:incoming_philo_slave_byteenable
	wire         mm_interconnect_0_philosopher_two_incoming_philo_slave_readdatavalid;  // philosopher_two:incoming_philo_slave_readdatavalid -> mm_interconnect_0:philosopher_two_incoming_philo_slave_readdatavalid
	wire         mm_interconnect_0_philosopher_two_incoming_philo_slave_write;          // mm_interconnect_0:philosopher_two_incoming_philo_slave_write -> philosopher_two:incoming_philo_slave_write
	wire  [31:0] mm_interconnect_0_philosopher_two_incoming_philo_slave_writedata;      // mm_interconnect_0:philosopher_two_incoming_philo_slave_writedata -> philosopher_two:incoming_philo_slave_writedata
	wire   [0:0] mm_interconnect_0_philosopher_two_incoming_philo_slave_burstcount;     // mm_interconnect_0:philosopher_two_incoming_philo_slave_burstcount -> philosopher_two:incoming_philo_slave_burstcount
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                         // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                           // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_s1_address;                            // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                         // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                              // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                          // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                              // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_timer_top_s1_chipselect;                             // mm_interconnect_0:timer_top_s1_chipselect -> timer_top:chipselect
	wire  [15:0] mm_interconnect_0_timer_top_s1_readdata;                               // timer_top:readdata -> mm_interconnect_0:timer_top_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_top_s1_address;                                // mm_interconnect_0:timer_top_s1_address -> timer_top:address
	wire         mm_interconnect_0_timer_top_s1_write;                                  // mm_interconnect_0:timer_top_s1_write -> timer_top:write_n
	wire  [15:0] mm_interconnect_0_timer_top_s1_writedata;                              // mm_interconnect_0:timer_top_s1_writedata -> timer_top:writedata
	wire         irq_mapper_receiver0_irq;                                              // timer_top:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                              // jtag_uart_top:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_top_irq_irq;                                                       // irq_mapper:sender_irq -> cpu_top:irq
	wire         rst_controller_reset_out_reset;                                        // rst_controller:reset_out -> [cpu_top:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_top_reset_reset_bridge_in_reset_reset, mm_interconnect_0:philosopher_zero_philosopher_clk_reset_in_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                                    // rst_controller:reset_req -> [cpu_top:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         philosopher_zero_cpu_jtag_debug_module_reset_reset;                    // philosopher_zero:cpu_jtag_debug_module_reset_reset -> [rst_controller:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in2]
	wire         philosopher_one_cpu_jtag_debug_module_reset_reset;                     // philosopher_one:cpu_jtag_debug_module_reset_reset -> [rst_controller:reset_in2, rst_controller_002:reset_in2, rst_controller_003:reset_in2, rst_controller_004:reset_in1]
	wire         philosopher_two_cpu_jtag_debug_module_reset_reset;                     // philosopher_two:cpu_jtag_debug_module_reset_reset -> [rst_controller:reset_in3, rst_controller_002:reset_in3, rst_controller_003:reset_in3, rst_controller_004:reset_in3]
	wire         cpu_top_debug_reset_request_reset;                                     // cpu_top:debug_reset_request -> [rst_controller:reset_in4, rst_controller_001:reset_in1, rst_controller_002:reset_in4, rst_controller_003:reset_in4, rst_controller_004:reset_in4]
	wire         rst_controller_001_reset_out_reset;                                    // rst_controller_001:reset_out -> [jtag_uart_top:rst_n, mm_interconnect_0:jtag_uart_top_reset_reset_bridge_in_reset_reset, timer_top:reset_n]
	wire         rst_controller_002_reset_out_reset;                                    // rst_controller_002:reset_out -> philosopher_one:philosopher_clk_reset_in_reset_n
	wire         rst_controller_003_reset_out_reset;                                    // rst_controller_003:reset_out -> philosopher_two:philosopher_clk_reset_in_reset_n
	wire         rst_controller_004_reset_out_reset;                                    // rst_controller_004:reset_out -> philosopher_zero:philosopher_clk_reset_in_reset_n

	multiprocessor_tutorial_main_system_cpu_top cpu_top (
		.clk                                 (clk_in_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (cpu_top_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_top_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_top_data_master_read),                              //                          .read
		.d_readdata                          (cpu_top_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_top_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_top_data_master_write),                             //                          .write
		.d_writedata                         (cpu_top_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_top_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_top_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_top_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_top_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_top_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_top_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_top_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_top_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_top_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_top_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_top_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_top_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_top_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_top_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_top_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	multiprocessor_tutorial_main_system_jtag_uart_top jtag_uart_top (
		.clk            (clk_in_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                       //               irq.irq
	);

	multiprocessor_tutorial_main_system_onchip_memory onchip_memory (
		.clk        (clk_in_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	multiprocessor_tutorial_main_system_philosopher_one philosopher_one (
		.cpu_jtag_debug_module_reset_reset   (philosopher_one_cpu_jtag_debug_module_reset_reset),                    // cpu_jtag_debug_module_reset.reset
		.incoming_philo_slave_waitrequest    (mm_interconnect_0_philosopher_one_incoming_philo_slave_waitrequest),   //        incoming_philo_slave.waitrequest
		.incoming_philo_slave_readdata       (mm_interconnect_0_philosopher_one_incoming_philo_slave_readdata),      //                            .readdata
		.incoming_philo_slave_readdatavalid  (mm_interconnect_0_philosopher_one_incoming_philo_slave_readdatavalid), //                            .readdatavalid
		.incoming_philo_slave_burstcount     (mm_interconnect_0_philosopher_one_incoming_philo_slave_burstcount),    //                            .burstcount
		.incoming_philo_slave_writedata      (mm_interconnect_0_philosopher_one_incoming_philo_slave_writedata),     //                            .writedata
		.incoming_philo_slave_address        (mm_interconnect_0_philosopher_one_incoming_philo_slave_address),       //                            .address
		.incoming_philo_slave_write          (mm_interconnect_0_philosopher_one_incoming_philo_slave_write),         //                            .write
		.incoming_philo_slave_read           (mm_interconnect_0_philosopher_one_incoming_philo_slave_read),          //                            .read
		.incoming_philo_slave_byteenable     (mm_interconnect_0_philosopher_one_incoming_philo_slave_byteenable),    //                            .byteenable
		.incoming_philo_slave_debugaccess    (mm_interconnect_0_philosopher_one_incoming_philo_slave_debugaccess),   //                            .debugaccess
		.outgoing_master_waitrequest         (philosopher_one_outgoing_master_waitrequest),                          //             outgoing_master.waitrequest
		.outgoing_master_readdata            (philosopher_one_outgoing_master_readdata),                             //                            .readdata
		.outgoing_master_readdatavalid       (philosopher_one_outgoing_master_readdatavalid),                        //                            .readdatavalid
		.outgoing_master_burstcount          (philosopher_one_outgoing_master_burstcount),                           //                            .burstcount
		.outgoing_master_writedata           (philosopher_one_outgoing_master_writedata),                            //                            .writedata
		.outgoing_master_address             (philosopher_one_outgoing_master_address),                              //                            .address
		.outgoing_master_write               (philosopher_one_outgoing_master_write),                                //                            .write
		.outgoing_master_read                (philosopher_one_outgoing_master_read),                                 //                            .read
		.outgoing_master_byteenable          (philosopher_one_outgoing_master_byteenable),                           //                            .byteenable
		.outgoing_master_debugaccess         (philosopher_one_outgoing_master_debugaccess),                          //                            .debugaccess
		.outgoing_philo_master_waitrequest   (philosopher_one_outgoing_philo_master_waitrequest),                    //       outgoing_philo_master.waitrequest
		.outgoing_philo_master_readdata      (philosopher_one_outgoing_philo_master_readdata),                       //                            .readdata
		.outgoing_philo_master_readdatavalid (philosopher_one_outgoing_philo_master_readdatavalid),                  //                            .readdatavalid
		.outgoing_philo_master_burstcount    (philosopher_one_outgoing_philo_master_burstcount),                     //                            .burstcount
		.outgoing_philo_master_writedata     (philosopher_one_outgoing_philo_master_writedata),                      //                            .writedata
		.outgoing_philo_master_address       (philosopher_one_outgoing_philo_master_address),                        //                            .address
		.outgoing_philo_master_write         (philosopher_one_outgoing_philo_master_write),                          //                            .write
		.outgoing_philo_master_read          (philosopher_one_outgoing_philo_master_read),                           //                            .read
		.outgoing_philo_master_byteenable    (philosopher_one_outgoing_philo_master_byteenable),                     //                            .byteenable
		.outgoing_philo_master_debugaccess   (philosopher_one_outgoing_philo_master_debugaccess),                    //                            .debugaccess
		.philosopher_clk_in_clk              (clk_in_clk),                                                           //          philosopher_clk_in.clk
		.philosopher_clk_reset_in_reset_n    (~rst_controller_002_reset_out_reset)                                   //    philosopher_clk_reset_in.reset_n
	);

	multiprocessor_tutorial_main_system_philosopher_two philosopher_two (
		.cpu_jtag_debug_module_reset_reset   (philosopher_two_cpu_jtag_debug_module_reset_reset),                    // cpu_jtag_debug_module_reset.reset
		.incoming_philo_slave_waitrequest    (mm_interconnect_0_philosopher_two_incoming_philo_slave_waitrequest),   //        incoming_philo_slave.waitrequest
		.incoming_philo_slave_readdata       (mm_interconnect_0_philosopher_two_incoming_philo_slave_readdata),      //                            .readdata
		.incoming_philo_slave_readdatavalid  (mm_interconnect_0_philosopher_two_incoming_philo_slave_readdatavalid), //                            .readdatavalid
		.incoming_philo_slave_burstcount     (mm_interconnect_0_philosopher_two_incoming_philo_slave_burstcount),    //                            .burstcount
		.incoming_philo_slave_writedata      (mm_interconnect_0_philosopher_two_incoming_philo_slave_writedata),     //                            .writedata
		.incoming_philo_slave_address        (mm_interconnect_0_philosopher_two_incoming_philo_slave_address),       //                            .address
		.incoming_philo_slave_write          (mm_interconnect_0_philosopher_two_incoming_philo_slave_write),         //                            .write
		.incoming_philo_slave_read           (mm_interconnect_0_philosopher_two_incoming_philo_slave_read),          //                            .read
		.incoming_philo_slave_byteenable     (mm_interconnect_0_philosopher_two_incoming_philo_slave_byteenable),    //                            .byteenable
		.incoming_philo_slave_debugaccess    (mm_interconnect_0_philosopher_two_incoming_philo_slave_debugaccess),   //                            .debugaccess
		.outgoing_master_waitrequest         (philosopher_two_outgoing_master_waitrequest),                          //             outgoing_master.waitrequest
		.outgoing_master_readdata            (philosopher_two_outgoing_master_readdata),                             //                            .readdata
		.outgoing_master_readdatavalid       (philosopher_two_outgoing_master_readdatavalid),                        //                            .readdatavalid
		.outgoing_master_burstcount          (philosopher_two_outgoing_master_burstcount),                           //                            .burstcount
		.outgoing_master_writedata           (philosopher_two_outgoing_master_writedata),                            //                            .writedata
		.outgoing_master_address             (philosopher_two_outgoing_master_address),                              //                            .address
		.outgoing_master_write               (philosopher_two_outgoing_master_write),                                //                            .write
		.outgoing_master_read                (philosopher_two_outgoing_master_read),                                 //                            .read
		.outgoing_master_byteenable          (philosopher_two_outgoing_master_byteenable),                           //                            .byteenable
		.outgoing_master_debugaccess         (philosopher_two_outgoing_master_debugaccess),                          //                            .debugaccess
		.outgoing_philo_master_waitrequest   (philosopher_two_outgoing_philo_master_waitrequest),                    //       outgoing_philo_master.waitrequest
		.outgoing_philo_master_readdata      (philosopher_two_outgoing_philo_master_readdata),                       //                            .readdata
		.outgoing_philo_master_readdatavalid (philosopher_two_outgoing_philo_master_readdatavalid),                  //                            .readdatavalid
		.outgoing_philo_master_burstcount    (philosopher_two_outgoing_philo_master_burstcount),                     //                            .burstcount
		.outgoing_philo_master_writedata     (philosopher_two_outgoing_philo_master_writedata),                      //                            .writedata
		.outgoing_philo_master_address       (philosopher_two_outgoing_philo_master_address),                        //                            .address
		.outgoing_philo_master_write         (philosopher_two_outgoing_philo_master_write),                          //                            .write
		.outgoing_philo_master_read          (philosopher_two_outgoing_philo_master_read),                           //                            .read
		.outgoing_philo_master_byteenable    (philosopher_two_outgoing_philo_master_byteenable),                     //                            .byteenable
		.outgoing_philo_master_debugaccess   (philosopher_two_outgoing_philo_master_debugaccess),                    //                            .debugaccess
		.philosopher_clk_in_clk              (clk_in_clk),                                                           //          philosopher_clk_in.clk
		.philosopher_clk_reset_in_reset_n    (~rst_controller_003_reset_out_reset)                                   //    philosopher_clk_reset_in.reset_n
	);

	multiprocessor_tutorial_main_system_philosopher_zero philosopher_zero (
		.cpu_jtag_debug_module_reset_reset   (philosopher_zero_cpu_jtag_debug_module_reset_reset),                    // cpu_jtag_debug_module_reset.reset
		.incoming_philo_slave_waitrequest    (mm_interconnect_0_philosopher_zero_incoming_philo_slave_waitrequest),   //        incoming_philo_slave.waitrequest
		.incoming_philo_slave_readdata       (mm_interconnect_0_philosopher_zero_incoming_philo_slave_readdata),      //                            .readdata
		.incoming_philo_slave_readdatavalid  (mm_interconnect_0_philosopher_zero_incoming_philo_slave_readdatavalid), //                            .readdatavalid
		.incoming_philo_slave_burstcount     (mm_interconnect_0_philosopher_zero_incoming_philo_slave_burstcount),    //                            .burstcount
		.incoming_philo_slave_writedata      (mm_interconnect_0_philosopher_zero_incoming_philo_slave_writedata),     //                            .writedata
		.incoming_philo_slave_address        (mm_interconnect_0_philosopher_zero_incoming_philo_slave_address),       //                            .address
		.incoming_philo_slave_write          (mm_interconnect_0_philosopher_zero_incoming_philo_slave_write),         //                            .write
		.incoming_philo_slave_read           (mm_interconnect_0_philosopher_zero_incoming_philo_slave_read),          //                            .read
		.incoming_philo_slave_byteenable     (mm_interconnect_0_philosopher_zero_incoming_philo_slave_byteenable),    //                            .byteenable
		.incoming_philo_slave_debugaccess    (mm_interconnect_0_philosopher_zero_incoming_philo_slave_debugaccess),   //                            .debugaccess
		.outgoing_master_waitrequest         (philosopher_zero_outgoing_master_waitrequest),                          //             outgoing_master.waitrequest
		.outgoing_master_readdata            (philosopher_zero_outgoing_master_readdata),                             //                            .readdata
		.outgoing_master_readdatavalid       (philosopher_zero_outgoing_master_readdatavalid),                        //                            .readdatavalid
		.outgoing_master_burstcount          (philosopher_zero_outgoing_master_burstcount),                           //                            .burstcount
		.outgoing_master_writedata           (philosopher_zero_outgoing_master_writedata),                            //                            .writedata
		.outgoing_master_address             (philosopher_zero_outgoing_master_address),                              //                            .address
		.outgoing_master_write               (philosopher_zero_outgoing_master_write),                                //                            .write
		.outgoing_master_read                (philosopher_zero_outgoing_master_read),                                 //                            .read
		.outgoing_master_byteenable          (philosopher_zero_outgoing_master_byteenable),                           //                            .byteenable
		.outgoing_master_debugaccess         (philosopher_zero_outgoing_master_debugaccess),                          //                            .debugaccess
		.outgoing_philo_master_waitrequest   (philosopher_zero_outgoing_philo_master_waitrequest),                    //       outgoing_philo_master.waitrequest
		.outgoing_philo_master_readdata      (philosopher_zero_outgoing_philo_master_readdata),                       //                            .readdata
		.outgoing_philo_master_readdatavalid (philosopher_zero_outgoing_philo_master_readdatavalid),                  //                            .readdatavalid
		.outgoing_philo_master_burstcount    (philosopher_zero_outgoing_philo_master_burstcount),                     //                            .burstcount
		.outgoing_philo_master_writedata     (philosopher_zero_outgoing_philo_master_writedata),                      //                            .writedata
		.outgoing_philo_master_address       (philosopher_zero_outgoing_philo_master_address),                        //                            .address
		.outgoing_philo_master_write         (philosopher_zero_outgoing_philo_master_write),                          //                            .write
		.outgoing_philo_master_read          (philosopher_zero_outgoing_philo_master_read),                           //                            .read
		.outgoing_philo_master_byteenable    (philosopher_zero_outgoing_philo_master_byteenable),                     //                            .byteenable
		.outgoing_philo_master_debugaccess   (philosopher_zero_outgoing_philo_master_debugaccess),                    //                            .debugaccess
		.philosopher_clk_in_clk              (clk_in_clk),                                                            //          philosopher_clk_in.clk
		.philosopher_clk_reset_in_reset_n    (~rst_controller_004_reset_out_reset)                                    //    philosopher_clk_reset_in.reset_n
	);

	multiprocessor_tutorial_main_system_sysid_qsys sysid_qsys (
		.clock    (clk_in_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	multiprocessor_tutorial_main_system_timer_top timer_top (
		.clk        (clk_in_clk),                                //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_top_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_top_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_top_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_top_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_top_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                   //   irq.irq
	);

	multiprocessor_tutorial_main_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                                           (clk_in_clk),                                                            //                                                         clk_clk.clk
		.cpu_top_reset_reset_bridge_in_reset_reset                             (rst_controller_reset_out_reset),                                        //                             cpu_top_reset_reset_bridge_in_reset.reset
		.jtag_uart_top_reset_reset_bridge_in_reset_reset                       (rst_controller_001_reset_out_reset),                                    //                       jtag_uart_top_reset_reset_bridge_in_reset.reset
		.philosopher_zero_philosopher_clk_reset_in_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                        // philosopher_zero_philosopher_clk_reset_in_reset_bridge_in_reset.reset
		.cpu_top_data_master_address                                           (cpu_top_data_master_address),                                           //                                             cpu_top_data_master.address
		.cpu_top_data_master_waitrequest                                       (cpu_top_data_master_waitrequest),                                       //                                                                .waitrequest
		.cpu_top_data_master_byteenable                                        (cpu_top_data_master_byteenable),                                        //                                                                .byteenable
		.cpu_top_data_master_read                                              (cpu_top_data_master_read),                                              //                                                                .read
		.cpu_top_data_master_readdata                                          (cpu_top_data_master_readdata),                                          //                                                                .readdata
		.cpu_top_data_master_write                                             (cpu_top_data_master_write),                                             //                                                                .write
		.cpu_top_data_master_writedata                                         (cpu_top_data_master_writedata),                                         //                                                                .writedata
		.cpu_top_data_master_debugaccess                                       (cpu_top_data_master_debugaccess),                                       //                                                                .debugaccess
		.cpu_top_instruction_master_address                                    (cpu_top_instruction_master_address),                                    //                                      cpu_top_instruction_master.address
		.cpu_top_instruction_master_waitrequest                                (cpu_top_instruction_master_waitrequest),                                //                                                                .waitrequest
		.cpu_top_instruction_master_read                                       (cpu_top_instruction_master_read),                                       //                                                                .read
		.cpu_top_instruction_master_readdata                                   (cpu_top_instruction_master_readdata),                                   //                                                                .readdata
		.philosopher_one_outgoing_master_address                               (philosopher_one_outgoing_master_address),                               //                                 philosopher_one_outgoing_master.address
		.philosopher_one_outgoing_master_waitrequest                           (philosopher_one_outgoing_master_waitrequest),                           //                                                                .waitrequest
		.philosopher_one_outgoing_master_burstcount                            (philosopher_one_outgoing_master_burstcount),                            //                                                                .burstcount
		.philosopher_one_outgoing_master_byteenable                            (philosopher_one_outgoing_master_byteenable),                            //                                                                .byteenable
		.philosopher_one_outgoing_master_read                                  (philosopher_one_outgoing_master_read),                                  //                                                                .read
		.philosopher_one_outgoing_master_readdata                              (philosopher_one_outgoing_master_readdata),                              //                                                                .readdata
		.philosopher_one_outgoing_master_readdatavalid                         (philosopher_one_outgoing_master_readdatavalid),                         //                                                                .readdatavalid
		.philosopher_one_outgoing_master_write                                 (philosopher_one_outgoing_master_write),                                 //                                                                .write
		.philosopher_one_outgoing_master_writedata                             (philosopher_one_outgoing_master_writedata),                             //                                                                .writedata
		.philosopher_one_outgoing_master_debugaccess                           (philosopher_one_outgoing_master_debugaccess),                           //                                                                .debugaccess
		.philosopher_one_outgoing_philo_master_address                         (philosopher_one_outgoing_philo_master_address),                         //                           philosopher_one_outgoing_philo_master.address
		.philosopher_one_outgoing_philo_master_waitrequest                     (philosopher_one_outgoing_philo_master_waitrequest),                     //                                                                .waitrequest
		.philosopher_one_outgoing_philo_master_burstcount                      (philosopher_one_outgoing_philo_master_burstcount),                      //                                                                .burstcount
		.philosopher_one_outgoing_philo_master_byteenable                      (philosopher_one_outgoing_philo_master_byteenable),                      //                                                                .byteenable
		.philosopher_one_outgoing_philo_master_read                            (philosopher_one_outgoing_philo_master_read),                            //                                                                .read
		.philosopher_one_outgoing_philo_master_readdata                        (philosopher_one_outgoing_philo_master_readdata),                        //                                                                .readdata
		.philosopher_one_outgoing_philo_master_readdatavalid                   (philosopher_one_outgoing_philo_master_readdatavalid),                   //                                                                .readdatavalid
		.philosopher_one_outgoing_philo_master_write                           (philosopher_one_outgoing_philo_master_write),                           //                                                                .write
		.philosopher_one_outgoing_philo_master_writedata                       (philosopher_one_outgoing_philo_master_writedata),                       //                                                                .writedata
		.philosopher_one_outgoing_philo_master_debugaccess                     (philosopher_one_outgoing_philo_master_debugaccess),                     //                                                                .debugaccess
		.philosopher_two_outgoing_master_address                               (philosopher_two_outgoing_master_address),                               //                                 philosopher_two_outgoing_master.address
		.philosopher_two_outgoing_master_waitrequest                           (philosopher_two_outgoing_master_waitrequest),                           //                                                                .waitrequest
		.philosopher_two_outgoing_master_burstcount                            (philosopher_two_outgoing_master_burstcount),                            //                                                                .burstcount
		.philosopher_two_outgoing_master_byteenable                            (philosopher_two_outgoing_master_byteenable),                            //                                                                .byteenable
		.philosopher_two_outgoing_master_read                                  (philosopher_two_outgoing_master_read),                                  //                                                                .read
		.philosopher_two_outgoing_master_readdata                              (philosopher_two_outgoing_master_readdata),                              //                                                                .readdata
		.philosopher_two_outgoing_master_readdatavalid                         (philosopher_two_outgoing_master_readdatavalid),                         //                                                                .readdatavalid
		.philosopher_two_outgoing_master_write                                 (philosopher_two_outgoing_master_write),                                 //                                                                .write
		.philosopher_two_outgoing_master_writedata                             (philosopher_two_outgoing_master_writedata),                             //                                                                .writedata
		.philosopher_two_outgoing_master_debugaccess                           (philosopher_two_outgoing_master_debugaccess),                           //                                                                .debugaccess
		.philosopher_two_outgoing_philo_master_address                         (philosopher_two_outgoing_philo_master_address),                         //                           philosopher_two_outgoing_philo_master.address
		.philosopher_two_outgoing_philo_master_waitrequest                     (philosopher_two_outgoing_philo_master_waitrequest),                     //                                                                .waitrequest
		.philosopher_two_outgoing_philo_master_burstcount                      (philosopher_two_outgoing_philo_master_burstcount),                      //                                                                .burstcount
		.philosopher_two_outgoing_philo_master_byteenable                      (philosopher_two_outgoing_philo_master_byteenable),                      //                                                                .byteenable
		.philosopher_two_outgoing_philo_master_read                            (philosopher_two_outgoing_philo_master_read),                            //                                                                .read
		.philosopher_two_outgoing_philo_master_readdata                        (philosopher_two_outgoing_philo_master_readdata),                        //                                                                .readdata
		.philosopher_two_outgoing_philo_master_readdatavalid                   (philosopher_two_outgoing_philo_master_readdatavalid),                   //                                                                .readdatavalid
		.philosopher_two_outgoing_philo_master_write                           (philosopher_two_outgoing_philo_master_write),                           //                                                                .write
		.philosopher_two_outgoing_philo_master_writedata                       (philosopher_two_outgoing_philo_master_writedata),                       //                                                                .writedata
		.philosopher_two_outgoing_philo_master_debugaccess                     (philosopher_two_outgoing_philo_master_debugaccess),                     //                                                                .debugaccess
		.philosopher_zero_outgoing_master_address                              (philosopher_zero_outgoing_master_address),                              //                                philosopher_zero_outgoing_master.address
		.philosopher_zero_outgoing_master_waitrequest                          (philosopher_zero_outgoing_master_waitrequest),                          //                                                                .waitrequest
		.philosopher_zero_outgoing_master_burstcount                           (philosopher_zero_outgoing_master_burstcount),                           //                                                                .burstcount
		.philosopher_zero_outgoing_master_byteenable                           (philosopher_zero_outgoing_master_byteenable),                           //                                                                .byteenable
		.philosopher_zero_outgoing_master_read                                 (philosopher_zero_outgoing_master_read),                                 //                                                                .read
		.philosopher_zero_outgoing_master_readdata                             (philosopher_zero_outgoing_master_readdata),                             //                                                                .readdata
		.philosopher_zero_outgoing_master_readdatavalid                        (philosopher_zero_outgoing_master_readdatavalid),                        //                                                                .readdatavalid
		.philosopher_zero_outgoing_master_write                                (philosopher_zero_outgoing_master_write),                                //                                                                .write
		.philosopher_zero_outgoing_master_writedata                            (philosopher_zero_outgoing_master_writedata),                            //                                                                .writedata
		.philosopher_zero_outgoing_master_debugaccess                          (philosopher_zero_outgoing_master_debugaccess),                          //                                                                .debugaccess
		.philosopher_zero_outgoing_philo_master_address                        (philosopher_zero_outgoing_philo_master_address),                        //                          philosopher_zero_outgoing_philo_master.address
		.philosopher_zero_outgoing_philo_master_waitrequest                    (philosopher_zero_outgoing_philo_master_waitrequest),                    //                                                                .waitrequest
		.philosopher_zero_outgoing_philo_master_burstcount                     (philosopher_zero_outgoing_philo_master_burstcount),                     //                                                                .burstcount
		.philosopher_zero_outgoing_philo_master_byteenable                     (philosopher_zero_outgoing_philo_master_byteenable),                     //                                                                .byteenable
		.philosopher_zero_outgoing_philo_master_read                           (philosopher_zero_outgoing_philo_master_read),                           //                                                                .read
		.philosopher_zero_outgoing_philo_master_readdata                       (philosopher_zero_outgoing_philo_master_readdata),                       //                                                                .readdata
		.philosopher_zero_outgoing_philo_master_readdatavalid                  (philosopher_zero_outgoing_philo_master_readdatavalid),                  //                                                                .readdatavalid
		.philosopher_zero_outgoing_philo_master_write                          (philosopher_zero_outgoing_philo_master_write),                          //                                                                .write
		.philosopher_zero_outgoing_philo_master_writedata                      (philosopher_zero_outgoing_philo_master_writedata),                      //                                                                .writedata
		.philosopher_zero_outgoing_philo_master_debugaccess                    (philosopher_zero_outgoing_philo_master_debugaccess),                    //                                                                .debugaccess
		.cpu_top_debug_mem_slave_address                                       (mm_interconnect_0_cpu_top_debug_mem_slave_address),                     //                                         cpu_top_debug_mem_slave.address
		.cpu_top_debug_mem_slave_write                                         (mm_interconnect_0_cpu_top_debug_mem_slave_write),                       //                                                                .write
		.cpu_top_debug_mem_slave_read                                          (mm_interconnect_0_cpu_top_debug_mem_slave_read),                        //                                                                .read
		.cpu_top_debug_mem_slave_readdata                                      (mm_interconnect_0_cpu_top_debug_mem_slave_readdata),                    //                                                                .readdata
		.cpu_top_debug_mem_slave_writedata                                     (mm_interconnect_0_cpu_top_debug_mem_slave_writedata),                   //                                                                .writedata
		.cpu_top_debug_mem_slave_byteenable                                    (mm_interconnect_0_cpu_top_debug_mem_slave_byteenable),                  //                                                                .byteenable
		.cpu_top_debug_mem_slave_waitrequest                                   (mm_interconnect_0_cpu_top_debug_mem_slave_waitrequest),                 //                                                                .waitrequest
		.cpu_top_debug_mem_slave_debugaccess                                   (mm_interconnect_0_cpu_top_debug_mem_slave_debugaccess),                 //                                                                .debugaccess
		.jtag_uart_top_avalon_jtag_slave_address                               (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_address),             //                                 jtag_uart_top_avalon_jtag_slave.address
		.jtag_uart_top_avalon_jtag_slave_write                                 (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_write),               //                                                                .write
		.jtag_uart_top_avalon_jtag_slave_read                                  (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_read),                //                                                                .read
		.jtag_uart_top_avalon_jtag_slave_readdata                              (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_readdata),            //                                                                .readdata
		.jtag_uart_top_avalon_jtag_slave_writedata                             (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_writedata),           //                                                                .writedata
		.jtag_uart_top_avalon_jtag_slave_waitrequest                           (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_waitrequest),         //                                                                .waitrequest
		.jtag_uart_top_avalon_jtag_slave_chipselect                            (mm_interconnect_0_jtag_uart_top_avalon_jtag_slave_chipselect),          //                                                                .chipselect
		.onchip_memory_s1_address                                              (mm_interconnect_0_onchip_memory_s1_address),                            //                                                onchip_memory_s1.address
		.onchip_memory_s1_write                                                (mm_interconnect_0_onchip_memory_s1_write),                              //                                                                .write
		.onchip_memory_s1_readdata                                             (mm_interconnect_0_onchip_memory_s1_readdata),                           //                                                                .readdata
		.onchip_memory_s1_writedata                                            (mm_interconnect_0_onchip_memory_s1_writedata),                          //                                                                .writedata
		.onchip_memory_s1_byteenable                                           (mm_interconnect_0_onchip_memory_s1_byteenable),                         //                                                                .byteenable
		.onchip_memory_s1_chipselect                                           (mm_interconnect_0_onchip_memory_s1_chipselect),                         //                                                                .chipselect
		.onchip_memory_s1_clken                                                (mm_interconnect_0_onchip_memory_s1_clken),                              //                                                                .clken
		.philosopher_one_incoming_philo_slave_address                          (mm_interconnect_0_philosopher_one_incoming_philo_slave_address),        //                            philosopher_one_incoming_philo_slave.address
		.philosopher_one_incoming_philo_slave_write                            (mm_interconnect_0_philosopher_one_incoming_philo_slave_write),          //                                                                .write
		.philosopher_one_incoming_philo_slave_read                             (mm_interconnect_0_philosopher_one_incoming_philo_slave_read),           //                                                                .read
		.philosopher_one_incoming_philo_slave_readdata                         (mm_interconnect_0_philosopher_one_incoming_philo_slave_readdata),       //                                                                .readdata
		.philosopher_one_incoming_philo_slave_writedata                        (mm_interconnect_0_philosopher_one_incoming_philo_slave_writedata),      //                                                                .writedata
		.philosopher_one_incoming_philo_slave_burstcount                       (mm_interconnect_0_philosopher_one_incoming_philo_slave_burstcount),     //                                                                .burstcount
		.philosopher_one_incoming_philo_slave_byteenable                       (mm_interconnect_0_philosopher_one_incoming_philo_slave_byteenable),     //                                                                .byteenable
		.philosopher_one_incoming_philo_slave_readdatavalid                    (mm_interconnect_0_philosopher_one_incoming_philo_slave_readdatavalid),  //                                                                .readdatavalid
		.philosopher_one_incoming_philo_slave_waitrequest                      (mm_interconnect_0_philosopher_one_incoming_philo_slave_waitrequest),    //                                                                .waitrequest
		.philosopher_one_incoming_philo_slave_debugaccess                      (mm_interconnect_0_philosopher_one_incoming_philo_slave_debugaccess),    //                                                                .debugaccess
		.philosopher_two_incoming_philo_slave_address                          (mm_interconnect_0_philosopher_two_incoming_philo_slave_address),        //                            philosopher_two_incoming_philo_slave.address
		.philosopher_two_incoming_philo_slave_write                            (mm_interconnect_0_philosopher_two_incoming_philo_slave_write),          //                                                                .write
		.philosopher_two_incoming_philo_slave_read                             (mm_interconnect_0_philosopher_two_incoming_philo_slave_read),           //                                                                .read
		.philosopher_two_incoming_philo_slave_readdata                         (mm_interconnect_0_philosopher_two_incoming_philo_slave_readdata),       //                                                                .readdata
		.philosopher_two_incoming_philo_slave_writedata                        (mm_interconnect_0_philosopher_two_incoming_philo_slave_writedata),      //                                                                .writedata
		.philosopher_two_incoming_philo_slave_burstcount                       (mm_interconnect_0_philosopher_two_incoming_philo_slave_burstcount),     //                                                                .burstcount
		.philosopher_two_incoming_philo_slave_byteenable                       (mm_interconnect_0_philosopher_two_incoming_philo_slave_byteenable),     //                                                                .byteenable
		.philosopher_two_incoming_philo_slave_readdatavalid                    (mm_interconnect_0_philosopher_two_incoming_philo_slave_readdatavalid),  //                                                                .readdatavalid
		.philosopher_two_incoming_philo_slave_waitrequest                      (mm_interconnect_0_philosopher_two_incoming_philo_slave_waitrequest),    //                                                                .waitrequest
		.philosopher_two_incoming_philo_slave_debugaccess                      (mm_interconnect_0_philosopher_two_incoming_philo_slave_debugaccess),    //                                                                .debugaccess
		.philosopher_zero_incoming_philo_slave_address                         (mm_interconnect_0_philosopher_zero_incoming_philo_slave_address),       //                           philosopher_zero_incoming_philo_slave.address
		.philosopher_zero_incoming_philo_slave_write                           (mm_interconnect_0_philosopher_zero_incoming_philo_slave_write),         //                                                                .write
		.philosopher_zero_incoming_philo_slave_read                            (mm_interconnect_0_philosopher_zero_incoming_philo_slave_read),          //                                                                .read
		.philosopher_zero_incoming_philo_slave_readdata                        (mm_interconnect_0_philosopher_zero_incoming_philo_slave_readdata),      //                                                                .readdata
		.philosopher_zero_incoming_philo_slave_writedata                       (mm_interconnect_0_philosopher_zero_incoming_philo_slave_writedata),     //                                                                .writedata
		.philosopher_zero_incoming_philo_slave_burstcount                      (mm_interconnect_0_philosopher_zero_incoming_philo_slave_burstcount),    //                                                                .burstcount
		.philosopher_zero_incoming_philo_slave_byteenable                      (mm_interconnect_0_philosopher_zero_incoming_philo_slave_byteenable),    //                                                                .byteenable
		.philosopher_zero_incoming_philo_slave_readdatavalid                   (mm_interconnect_0_philosopher_zero_incoming_philo_slave_readdatavalid), //                                                                .readdatavalid
		.philosopher_zero_incoming_philo_slave_waitrequest                     (mm_interconnect_0_philosopher_zero_incoming_philo_slave_waitrequest),   //                                                                .waitrequest
		.philosopher_zero_incoming_philo_slave_debugaccess                     (mm_interconnect_0_philosopher_zero_incoming_philo_slave_debugaccess),   //                                                                .debugaccess
		.sysid_qsys_control_slave_address                                      (mm_interconnect_0_sysid_qsys_control_slave_address),                    //                                        sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                     (mm_interconnect_0_sysid_qsys_control_slave_readdata),                   //                                                                .readdata
		.timer_top_s1_address                                                  (mm_interconnect_0_timer_top_s1_address),                                //                                                    timer_top_s1.address
		.timer_top_s1_write                                                    (mm_interconnect_0_timer_top_s1_write),                                  //                                                                .write
		.timer_top_s1_readdata                                                 (mm_interconnect_0_timer_top_s1_readdata),                               //                                                                .readdata
		.timer_top_s1_writedata                                                (mm_interconnect_0_timer_top_s1_writedata),                              //                                                                .writedata
		.timer_top_s1_chipselect                                               (mm_interconnect_0_timer_top_s1_chipselect)                              //                                                                .chipselect
	);

	multiprocessor_tutorial_main_system_irq_mapper irq_mapper (
		.clk           (clk_in_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_top_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (5),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clk_clk_in_reset_reset_n),                          // reset_in0.reset
		.reset_in1      (philosopher_zero_cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (philosopher_one_cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.reset_in3      (philosopher_two_cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.reset_in4      (cpu_top_debug_reset_request_reset),                  // reset_in4.reset
		.clk            (clk_in_clk),                                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),                 //          .reset_req
		.reset_req_in0  (1'b0),                                               // (terminated)
		.reset_req_in1  (1'b0),                                               // (terminated)
		.reset_req_in2  (1'b0),                                               // (terminated)
		.reset_req_in3  (1'b0),                                               // (terminated)
		.reset_req_in4  (1'b0),                                               // (terminated)
		.reset_in5      (1'b0),                                               // (terminated)
		.reset_req_in5  (1'b0),                                               // (terminated)
		.reset_in6      (1'b0),                                               // (terminated)
		.reset_req_in6  (1'b0),                                               // (terminated)
		.reset_in7      (1'b0),                                               // (terminated)
		.reset_req_in7  (1'b0),                                               // (terminated)
		.reset_in8      (1'b0),                                               // (terminated)
		.reset_req_in8  (1'b0),                                               // (terminated)
		.reset_in9      (1'b0),                                               // (terminated)
		.reset_req_in9  (1'b0),                                               // (terminated)
		.reset_in10     (1'b0),                                               // (terminated)
		.reset_req_in10 (1'b0),                                               // (terminated)
		.reset_in11     (1'b0),                                               // (terminated)
		.reset_req_in11 (1'b0),                                               // (terminated)
		.reset_in12     (1'b0),                                               // (terminated)
		.reset_req_in12 (1'b0),                                               // (terminated)
		.reset_in13     (1'b0),                                               // (terminated)
		.reset_req_in13 (1'b0),                                               // (terminated)
		.reset_in14     (1'b0),                                               // (terminated)
		.reset_req_in14 (1'b0),                                               // (terminated)
		.reset_in15     (1'b0),                                               // (terminated)
		.reset_req_in15 (1'b0)                                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~clk_clk_in_reset_reset_n),          // reset_in0.reset
		.reset_in1      (cpu_top_debug_reset_request_reset),  // reset_in1.reset
		.clk            (clk_in_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (5),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~clk_clk_in_reset_reset_n),                          // reset_in0.reset
		.reset_in1      (philosopher_zero_cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (philosopher_one_cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.reset_in3      (philosopher_two_cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.reset_in4      (cpu_top_debug_reset_request_reset),                  // reset_in4.reset
		.clk            (),                                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),                 // reset_out.reset
		.reset_req      (),                                                   // (terminated)
		.reset_req_in0  (1'b0),                                               // (terminated)
		.reset_req_in1  (1'b0),                                               // (terminated)
		.reset_req_in2  (1'b0),                                               // (terminated)
		.reset_req_in3  (1'b0),                                               // (terminated)
		.reset_req_in4  (1'b0),                                               // (terminated)
		.reset_in5      (1'b0),                                               // (terminated)
		.reset_req_in5  (1'b0),                                               // (terminated)
		.reset_in6      (1'b0),                                               // (terminated)
		.reset_req_in6  (1'b0),                                               // (terminated)
		.reset_in7      (1'b0),                                               // (terminated)
		.reset_req_in7  (1'b0),                                               // (terminated)
		.reset_in8      (1'b0),                                               // (terminated)
		.reset_req_in8  (1'b0),                                               // (terminated)
		.reset_in9      (1'b0),                                               // (terminated)
		.reset_req_in9  (1'b0),                                               // (terminated)
		.reset_in10     (1'b0),                                               // (terminated)
		.reset_req_in10 (1'b0),                                               // (terminated)
		.reset_in11     (1'b0),                                               // (terminated)
		.reset_req_in11 (1'b0),                                               // (terminated)
		.reset_in12     (1'b0),                                               // (terminated)
		.reset_req_in12 (1'b0),                                               // (terminated)
		.reset_in13     (1'b0),                                               // (terminated)
		.reset_req_in13 (1'b0),                                               // (terminated)
		.reset_in14     (1'b0),                                               // (terminated)
		.reset_req_in14 (1'b0),                                               // (terminated)
		.reset_in15     (1'b0),                                               // (terminated)
		.reset_req_in15 (1'b0)                                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (5),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~clk_clk_in_reset_reset_n),                          // reset_in0.reset
		.reset_in1      (philosopher_zero_cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (philosopher_one_cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.reset_in3      (philosopher_two_cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.reset_in4      (cpu_top_debug_reset_request_reset),                  // reset_in4.reset
		.clk            (),                                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),                 // reset_out.reset
		.reset_req      (),                                                   // (terminated)
		.reset_req_in0  (1'b0),                                               // (terminated)
		.reset_req_in1  (1'b0),                                               // (terminated)
		.reset_req_in2  (1'b0),                                               // (terminated)
		.reset_req_in3  (1'b0),                                               // (terminated)
		.reset_req_in4  (1'b0),                                               // (terminated)
		.reset_in5      (1'b0),                                               // (terminated)
		.reset_req_in5  (1'b0),                                               // (terminated)
		.reset_in6      (1'b0),                                               // (terminated)
		.reset_req_in6  (1'b0),                                               // (terminated)
		.reset_in7      (1'b0),                                               // (terminated)
		.reset_req_in7  (1'b0),                                               // (terminated)
		.reset_in8      (1'b0),                                               // (terminated)
		.reset_req_in8  (1'b0),                                               // (terminated)
		.reset_in9      (1'b0),                                               // (terminated)
		.reset_req_in9  (1'b0),                                               // (terminated)
		.reset_in10     (1'b0),                                               // (terminated)
		.reset_req_in10 (1'b0),                                               // (terminated)
		.reset_in11     (1'b0),                                               // (terminated)
		.reset_req_in11 (1'b0),                                               // (terminated)
		.reset_in12     (1'b0),                                               // (terminated)
		.reset_req_in12 (1'b0),                                               // (terminated)
		.reset_in13     (1'b0),                                               // (terminated)
		.reset_req_in13 (1'b0),                                               // (terminated)
		.reset_in14     (1'b0),                                               // (terminated)
		.reset_req_in14 (1'b0),                                               // (terminated)
		.reset_in15     (1'b0),                                               // (terminated)
		.reset_req_in15 (1'b0)                                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (5),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~clk_clk_in_reset_reset_n),                          // reset_in0.reset
		.reset_in1      (philosopher_one_cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.reset_in2      (philosopher_zero_cpu_jtag_debug_module_reset_reset), // reset_in2.reset
		.reset_in3      (philosopher_two_cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.reset_in4      (cpu_top_debug_reset_request_reset),                  // reset_in4.reset
		.clk            (),                                                   //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),                 // reset_out.reset
		.reset_req      (),                                                   // (terminated)
		.reset_req_in0  (1'b0),                                               // (terminated)
		.reset_req_in1  (1'b0),                                               // (terminated)
		.reset_req_in2  (1'b0),                                               // (terminated)
		.reset_req_in3  (1'b0),                                               // (terminated)
		.reset_req_in4  (1'b0),                                               // (terminated)
		.reset_in5      (1'b0),                                               // (terminated)
		.reset_req_in5  (1'b0),                                               // (terminated)
		.reset_in6      (1'b0),                                               // (terminated)
		.reset_req_in6  (1'b0),                                               // (terminated)
		.reset_in7      (1'b0),                                               // (terminated)
		.reset_req_in7  (1'b0),                                               // (terminated)
		.reset_in8      (1'b0),                                               // (terminated)
		.reset_req_in8  (1'b0),                                               // (terminated)
		.reset_in9      (1'b0),                                               // (terminated)
		.reset_req_in9  (1'b0),                                               // (terminated)
		.reset_in10     (1'b0),                                               // (terminated)
		.reset_req_in10 (1'b0),                                               // (terminated)
		.reset_in11     (1'b0),                                               // (terminated)
		.reset_req_in11 (1'b0),                                               // (terminated)
		.reset_in12     (1'b0),                                               // (terminated)
		.reset_req_in12 (1'b0),                                               // (terminated)
		.reset_in13     (1'b0),                                               // (terminated)
		.reset_req_in13 (1'b0),                                               // (terminated)
		.reset_in14     (1'b0),                                               // (terminated)
		.reset_req_in14 (1'b0),                                               // (terminated)
		.reset_in15     (1'b0),                                               // (terminated)
		.reset_req_in15 (1'b0)                                                // (terminated)
	);

endmodule
